module mul_signed (a,b,z); // 16x16 signed multiplier
	input [15:0] a, b; // a, b
	output [31:0] z; // z = a * b
	
	wire [15:0] ab0 = a & {16{b[0]}}; // a or 0 for b[0]
	wire [15:0] ab1 = a & {16{b[1]}}; // a or 0 for b[1]
	wire [15:0] ab2 = a & {16{b[2]}}; // a or 0 for b[2]
	wire [15:0] ab3 = a & {16{b[3]}}; // a or 0 for b[3]
	wire [15:0] ab4 = a & {16{b[4]}}; // a or 0 for b[4]
	wire [15:0] ab5 = a & {16{b[5]}}; // a or 0 for b[5]
	wire [15:0] ab6 = a & {16{b[6]}}; // a or 0 for b[6]
	wire [15:0] ab7 = a & {16{b[7]}}; // a or 0 for b[7]
	wire [15:0] ab8 = a & {16{b[8]}}; // a or 0 for b[0]
	wire [15:0] ab9 = a & {16{b[9]}}; // a or 0 for b[1]
	wire [15:0] ab10 = a & {16{b[10]}}; // a or 0 for b[2]
	wire [15:0] ab11 = a & {16{b[11]}}; // a or 0 for b[3]
	wire [15:0] ab12 = a & {16{b[12]}}; // a or 0 for b[4]
	wire [15:0] ab13 = a & {16{b[13]}}; // a or 0 for b[5]
	wire [15:0] ab14 = a & {16{b[14]}}; // a or 0 for b[6]
	wire [15:0] ab15 = a & {16{b[15]}}; // a or 0 for b[7]
	
	assign z = (({16'b1, ~ab0[15],   ab0[14:0]}               +   // << 0, + 1 in bit 16
					 {15'b0, ~ab1[15],   ab1[14:0],  1'b0})   +   // << 1
					({14'b0, ~ab2[15],   ab2[14:0],  2'b0}    +   // << 2
					 {13'b0, ~ab3[15],   ab3[14:0],  3'b0}))  +   // << 3
					(({12'b0,~ab4[15],   ab4[14:0],  4'b0}    +   // << 4
					 {11'b0, ~ab5[15],   ab5[14:0],  5'b0})   +   // << 5
					({10'b0, ~ab6[15],   ab6[14:0],  6'b0}    +   // << 6
					 {9'b0,  ~ab7[15],   ab7[14:0],  7'b0}))  +   // << 7
				  (({8'b0,  ~ab8[15],   ab8[14:0],  8'b0}     +   // << 8
					 {7'b0,  ~ab9[15],   ab9[14:0],  9'b0})   +   // << 9
					({6'b0,  ~ab10[15],  ab10[14:0],  10'b0}  +   // << 10
					 {5'b0,  ~ab11[15],  ab11[14:0],  11'b0}))+   // << 11
				  (({4'b0,  ~ab12[15],  ab12[14:0],  12'b0}   +   // << 12
					 {3'b0,  ~ab13[15],  ab13[14:0],  13'b0}) +   // << 13
					({2'b0,  ~ab14[15],  ab14[14:0],  14'b0}  +   // << 14
					 {1'b1,   ab15[15], ~ab15[14:0],  15'b0}));   // << 15, + 1 in bit 31
endmodule