module poolbanks(clk, rst, wren, rden, address, address2, datain, dataout);
input clk, rst;
reg [15:0] bank1 [0:111*111-1];
reg [15:0] bank2 [0:111*111-1];
reg [15:0] bank3 [0:111*111-1];
reg [15:0] bank4 [0:111*111-1];
reg [15:0] bank5 [0:111*111-1];
reg [15:0] bank6 [0:111*111-1];
reg [15:0] bank7 [0:111*111-1];
reg [15:0] bank8 [0:111*111-1];
reg [15:0] bank9 [0:111*111-1];
reg [15:0] bank10 [0:111*111-1];
reg [15:0] bank11 [0:111*111-1];
reg [15:0] bank12 [0:111*111-1];
reg [15:0] bank13 [0:111*111-1];
reg [15:0] bank14 [0:111*111-1];
reg [15:0] bank15 [0:111*111-1];
reg [15:0] bank16 [0:111*111-1];
reg [15:0] bank17 [0:111*111-1];
reg [15:0] bank18 [0:111*111-1];
reg [15:0] bank19 [0:111*111-1];
reg [15:0] bank20 [0:111*111-1];
reg [15:0] bank21 [0:111*111-1];
reg [15:0] bank22 [0:111*111-1];
reg [15:0] bank23 [0:111*111-1];
reg [15:0] bank24 [0:111*111-1];
reg [15:0] bank25 [0:111*111-1];
reg [15:0] bank26 [0:111*111-1];
reg [15:0] bank27 [0:111*111-1];
reg [15:0] bank28 [0:111*111-1];
reg [15:0] bank29 [0:111*111-1];
reg [15:0] bank30 [0:111*111-1];
reg [15:0] bank31 [0:111*111-1];
reg [15:0] bank32 [0:111*111-1];
reg [15:0] bank33 [0:111*111-1];
reg [15:0] bank34 [0:111*111-1];
reg [15:0] bank35 [0:111*111-1];
reg [15:0] bank36 [0:111*111-1];
reg [15:0] bank37 [0:111*111-1];
reg [15:0] bank38 [0:111*111-1];
reg [15:0] bank39 [0:111*111-1];
reg [15:0] bank40 [0:111*111-1];
reg [15:0] bank41 [0:111*111-1];
reg [15:0] bank42 [0:111*111-1];
reg [15:0] bank43 [0:111*111-1];
reg [15:0] bank44 [0:111*111-1];
reg [15:0] bank45 [0:111*111-1];
reg [15:0] bank46 [0:111*111-1];
reg [15:0] bank47 [0:111*111-1];
reg [15:0] bank48 [0:111*111-1];
reg [15:0] bank49 [0:111*111-1];
reg [15:0] bank50 [0:111*111-1];
reg [15:0] bank51 [0:111*111-1];
reg [15:0] bank52 [0:111*111-1];
reg [15:0] bank53 [0:111*111-1];
reg [15:0] bank54 [0:111*111-1];
reg [15:0] bank55 [0:111*111-1];
reg [15:0] bank56 [0:111*111-1];
reg [15:0] bank57 [0:111*111-1];
reg [15:0] bank58 [0:111*111-1];
reg [15:0] bank59 [0:111*111-1];
reg [15:0] bank60 [0:111*111-1];
reg [15:0] bank61 [0:111*111-1];
reg [15:0] bank62 [0:111*111-1];
reg [15:0] bank63 [0:111*111-1];
reg [15:0] bank64 [0:111*111-1];
reg [15:0] bank65 [0:111*111-1];
reg [15:0] bank66 [0:111*111-1];
reg [15:0] bank67 [0:111*111-1];
reg [15:0] bank68 [0:111*111-1];
reg [15:0] bank69 [0:111*111-1];
reg [15:0] bank70 [0:111*111-1];
reg [15:0] bank71 [0:111*111-1];
reg [15:0] bank72 [0:111*111-1];
reg [15:0] bank73 [0:111*111-1];
reg [15:0] bank74 [0:111*111-1];
reg [15:0] bank75 [0:111*111-1];
reg [15:0] bank76 [0:111*111-1];
reg [15:0] bank77 [0:111*111-1];
reg [15:0] bank78 [0:111*111-1];
reg [15:0] bank79 [0:111*111-1];
reg [15:0] bank80 [0:111*111-1];
reg [15:0] bank81 [0:111*111-1];
reg [15:0] bank82 [0:111*111-1];
reg [15:0] bank83 [0:111*111-1];
reg [15:0] bank84 [0:111*111-1];
reg [15:0] bank85 [0:111*111-1];
reg [15:0] bank86 [0:111*111-1];
reg [15:0] bank87 [0:111*111-1];
reg [15:0] bank88 [0:111*111-1];
reg [15:0] bank89 [0:111*111-1];
reg [15:0] bank90 [0:111*111-1];
reg [15:0] bank91 [0:111*111-1];
reg [15:0] bank92 [0:111*111-1];
reg [15:0] bank93 [0:111*111-1];
reg [15:0] bank94 [0:111*111-1];
reg [15:0] bank95 [0:111*111-1];
reg [15:0] bank96 [0:111*111-1];
reg [15:0] bank97 [0:111*111-1];
reg [15:0] bank98 [0:111*111-1];
reg [15:0] bank99 [0:111*111-1];
reg [15:0] bank100 [0:111*111-1];
reg [15:0] bank101 [0:111*111-1];
reg [15:0] bank102 [0:111*111-1];
reg [15:0] bank103 [0:111*111-1];
reg [15:0] bank104 [0:111*111-1];
reg [15:0] bank105 [0:111*111-1];
reg [15:0] bank106 [0:111*111-1];
reg [15:0] bank107 [0:111*111-1];
reg [15:0] bank108 [0:111*111-1];
reg [15:0] bank109 [0:111*111-1];
reg [15:0] bank110 [0:111*111-1];
reg [15:0] bank111 [0:111*111-1];
reg [15:0] bank112 [0:111*111-1];
reg [15:0] bank113 [0:111*111-1];
reg [15:0] bank114 [0:111*111-1];
reg [15:0] bank115 [0:111*111-1];
reg [15:0] bank116 [0:111*111-1];
reg [15:0] bank117 [0:111*111-1];
reg [15:0] bank118 [0:111*111-1];
reg [15:0] bank119 [0:111*111-1];
reg [15:0] bank120 [0:111*111-1];
reg [15:0] bank121 [0:111*111-1];
reg [15:0] bank122 [0:111*111-1];
reg [15:0] bank123 [0:111*111-1];
reg [15:0] bank124 [0:111*111-1];
reg [15:0] bank125 [0:111*111-1];
reg [15:0] bank126 [0:111*111-1];
reg [15:0] bank127 [0:111*111-1];
reg [15:0] bank128 [0:111*111-1];
reg [15:0] bank129 [0:111*111-1];
reg [15:0] bank130 [0:111*111-1];
reg [15:0] bank131 [0:111*111-1];
reg [15:0] bank132 [0:111*111-1];
reg [15:0] bank133 [0:111*111-1];
reg [15:0] bank134 [0:111*111-1];
reg [15:0] bank135 [0:111*111-1];
reg [15:0] bank136 [0:111*111-1];
reg [15:0] bank137 [0:111*111-1];
reg [15:0] bank138 [0:111*111-1];
reg [15:0] bank139 [0:111*111-1];
reg [15:0] bank140 [0:111*111-1];
reg [15:0] bank141 [0:111*111-1];
reg [15:0] bank142 [0:111*111-1];
reg [15:0] bank143 [0:111*111-1];
reg [15:0] bank144 [0:111*111-1];
reg [15:0] bank145 [0:111*111-1];
reg [15:0] bank146 [0:111*111-1];
reg [15:0] bank147 [0:111*111-1];
reg [15:0] bank148 [0:111*111-1];
reg [15:0] bank149 [0:111*111-1];
reg [15:0] bank150 [0:111*111-1];
reg [15:0] bank151 [0:111*111-1];
reg [15:0] bank152 [0:111*111-1];
reg [15:0] bank153 [0:111*111-1];
reg [15:0] bank154 [0:111*111-1];
reg [15:0] bank155 [0:111*111-1];
reg [15:0] bank156 [0:111*111-1];
reg [15:0] bank157 [0:111*111-1];
reg [15:0] bank158 [0:111*111-1];
reg [15:0] bank159 [0:111*111-1];
reg [15:0] bank160 [0:111*111-1];
reg [15:0] bank161 [0:111*111-1];
reg [15:0] bank162 [0:111*111-1];
reg [15:0] bank163 [0:111*111-1];
reg [15:0] bank164 [0:111*111-1];
reg [15:0] bank165 [0:111*111-1];
reg [15:0] bank166 [0:111*111-1];
reg [15:0] bank167 [0:111*111-1];
reg [15:0] bank168 [0:111*111-1];
reg [15:0] bank169 [0:111*111-1];
reg [15:0] bank170 [0:111*111-1];
reg [15:0] bank171 [0:111*111-1];
reg [15:0] bank172 [0:111*111-1];
reg [15:0] bank173 [0:111*111-1];
reg [15:0] bank174 [0:111*111-1];
reg [15:0] bank175 [0:111*111-1];
reg [15:0] bank176 [0:111*111-1];
reg [15:0] bank177 [0:111*111-1];
reg [15:0] bank178 [0:111*111-1];
reg [15:0] bank179 [0:111*111-1];
reg [15:0] bank180 [0:111*111-1];
reg [15:0] bank181 [0:111*111-1];
reg [15:0] bank182 [0:111*111-1];
reg [15:0] bank183 [0:111*111-1];
reg [15:0] bank184 [0:111*111-1];
reg [15:0] bank185 [0:111*111-1];
reg [15:0] bank186 [0:111*111-1];
reg [15:0] bank187 [0:111*111-1];
reg [15:0] bank188 [0:111*111-1];
reg [15:0] bank189 [0:111*111-1];
reg [15:0] bank190 [0:111*111-1];
reg [15:0] bank191 [0:111*111-1];
reg [15:0] bank192 [0:111*111-1];
reg [15:0] bank193 [0:111*111-1];
reg [15:0] bank194 [0:111*111-1];
reg [15:0] bank195 [0:111*111-1];
reg [15:0] bank196 [0:111*111-1];
reg [15:0] bank197 [0:111*111-1];
reg [15:0] bank198 [0:111*111-1];
reg [15:0] bank199 [0:111*111-1];
reg [15:0] bank200 [0:111*111-1];
reg [15:0] bank201 [0:111*111-1];
reg [15:0] bank202 [0:111*111-1];
reg [15:0] bank203 [0:111*111-1];
reg [15:0] bank204 [0:111*111-1];
reg [15:0] bank205 [0:111*111-1];
reg [15:0] bank206 [0:111*111-1];
reg [15:0] bank207 [0:111*111-1];
reg [15:0] bank208 [0:111*111-1];
reg [15:0] bank209 [0:111*111-1];
reg [15:0] bank210 [0:111*111-1];
reg [15:0] bank211 [0:111*111-1];
reg [15:0] bank212 [0:111*111-1];
reg [15:0] bank213 [0:111*111-1];
reg [15:0] bank214 [0:111*111-1];
reg [15:0] bank215 [0:111*111-1];
reg [15:0] bank216 [0:111*111-1];
reg [15:0] bank217 [0:111*111-1];
reg [15:0] bank218 [0:111*111-1];
reg [15:0] bank219 [0:111*111-1];
reg [15:0] bank220 [0:111*111-1];
reg [15:0] bank221 [0:111*111-1];
reg [15:0] bank222 [0:111*111-1];
reg [15:0] bank223 [0:111*111-1];
reg [15:0] bank224 [0:111*111-1];
reg [15:0] bank225 [0:111*111-1];
reg [15:0] bank226 [0:111*111-1];
reg [15:0] bank227 [0:111*111-1];
reg [15:0] bank228 [0:111*111-1];
reg [15:0] bank229 [0:111*111-1];
reg [15:0] bank230 [0:111*111-1];
reg [15:0] bank231 [0:111*111-1];
reg [15:0] bank232 [0:111*111-1];
reg [15:0] bank233 [0:111*111-1];
reg [15:0] bank234 [0:111*111-1];
reg [15:0] bank235 [0:111*111-1];
reg [15:0] bank236 [0:111*111-1];
reg [15:0] bank237 [0:111*111-1];
reg [15:0] bank238 [0:111*111-1];
reg [15:0] bank239 [0:111*111-1];
reg [15:0] bank240 [0:111*111-1];
reg [15:0] bank241 [0:111*111-1];
reg [15:0] bank242 [0:111*111-1];
reg [15:0] bank243 [0:111*111-1];
reg [15:0] bank244 [0:111*111-1];
reg [15:0] bank245 [0:111*111-1];
reg [15:0] bank246 [0:111*111-1];
reg [15:0] bank247 [0:111*111-1];
reg [15:0] bank248 [0:111*111-1];
reg [15:0] bank249 [0:111*111-1];
reg [15:0] bank250 [0:111*111-1];
reg [15:0] bank251 [0:111*111-1];
reg [15:0] bank252 [0:111*111-1];
reg [15:0] bank253 [0:111*111-1];
reg [15:0] bank254 [0:111*111-1];
reg [15:0] bank255 [0:111*111-1];
reg [15:0] bank256 [0:111*111-1];
input rden;
input wren;
input [32-1:0] address;
input [32-1:0] address2;
input [16*256-1:0] datain;
reg [15:0] datainmem[0:255];
output reg [16*256-1:0] dataout;
reg [15:0] dataoutmem[0:255];
integer i;
always @(*)
begin
for (i=0; i<256; i=i+1)
    datainmem[i]<=datain[i*16+:16];
end

always @(posedge clk)
begin
    if(rst)
        for (i=0; i<256;i=i+1) begin
            bank1[i] <= 16'd0;
            bank2[i] <= 16'd0;
            bank3[i] <= 16'd0;
            bank4[i] <= 16'd0;
            bank5[i] <= 16'd0;
            bank6[i] <= 16'd0;
            bank7[i] <= 16'd0;
            bank8[i] <= 16'd0;
            bank9[i] <= 16'd0;
            bank10[i] <= 16'd0;
            bank11[i] <= 16'd0;
            bank12[i] <= 16'd0;
            bank13[i] <= 16'd0;
            bank14[i] <= 16'd0;
            bank15[i] <= 16'd0;
            bank16[i] <= 16'd0;
            bank17[i] <= 16'd0;
            bank18[i] <= 16'd0;
            bank19[i] <= 16'd0;
            bank20[i] <= 16'd0;
            bank21[i] <= 16'd0;
            bank22[i] <= 16'd0;
            bank23[i] <= 16'd0;
            bank24[i] <= 16'd0;
            bank25[i] <= 16'd0;
            bank26[i] <= 16'd0;
            bank27[i] <= 16'd0;
            bank28[i] <= 16'd0;
            bank29[i] <= 16'd0;
            bank30[i] <= 16'd0;
            bank31[i] <= 16'd0;
            bank32[i] <= 16'd0;
            bank33[i] <= 16'd0;
            bank34[i] <= 16'd0;
            bank35[i] <= 16'd0;
            bank36[i] <= 16'd0;
            bank37[i] <= 16'd0;
            bank38[i] <= 16'd0;
            bank39[i] <= 16'd0;
            bank40[i] <= 16'd0;
            bank41[i] <= 16'd0;
            bank42[i] <= 16'd0;
            bank43[i] <= 16'd0;
            bank44[i] <= 16'd0;
            bank45[i] <= 16'd0;
            bank46[i] <= 16'd0;
            bank47[i] <= 16'd0;
            bank48[i] <= 16'd0;
            bank49[i] <= 16'd0;
            bank50[i] <= 16'd0;
            bank51[i] <= 16'd0;
            bank52[i] <= 16'd0;
            bank53[i] <= 16'd0;
            bank54[i] <= 16'd0;
            bank55[i] <= 16'd0;
            bank56[i] <= 16'd0;
            bank57[i] <= 16'd0;
            bank58[i] <= 16'd0;
            bank59[i] <= 16'd0;
            bank60[i] <= 16'd0;
            bank61[i] <= 16'd0;
            bank62[i] <= 16'd0;
            bank63[i] <= 16'd0;
            bank64[i] <= 16'd0;
            bank65[i] <= 16'd0;
            bank66[i] <= 16'd0;
            bank67[i] <= 16'd0;
            bank68[i] <= 16'd0;
            bank69[i] <= 16'd0;
            bank70[i] <= 16'd0;
            bank71[i] <= 16'd0;
            bank72[i] <= 16'd0;
            bank73[i] <= 16'd0;
            bank74[i] <= 16'd0;
            bank75[i] <= 16'd0;
            bank76[i] <= 16'd0;
            bank77[i] <= 16'd0;
            bank78[i] <= 16'd0;
            bank79[i] <= 16'd0;
            bank80[i] <= 16'd0;
            bank81[i] <= 16'd0;
            bank82[i] <= 16'd0;
            bank83[i] <= 16'd0;
            bank84[i] <= 16'd0;
            bank85[i] <= 16'd0;
            bank86[i] <= 16'd0;
            bank87[i] <= 16'd0;
            bank88[i] <= 16'd0;
            bank89[i] <= 16'd0;
            bank90[i] <= 16'd0;
            bank91[i] <= 16'd0;
            bank92[i] <= 16'd0;
            bank93[i] <= 16'd0;
            bank94[i] <= 16'd0;
            bank95[i] <= 16'd0;
            bank96[i] <= 16'd0;
            bank97[i] <= 16'd0;
            bank98[i] <= 16'd0;
            bank99[i] <= 16'd0;
            bank100[i] <= 16'd0;
            bank101[i] <= 16'd0;
            bank102[i] <= 16'd0;
            bank103[i] <= 16'd0;
            bank104[i] <= 16'd0;
            bank105[i] <= 16'd0;
            bank106[i] <= 16'd0;
            bank107[i] <= 16'd0;
            bank108[i] <= 16'd0;
            bank109[i] <= 16'd0;
            bank110[i] <= 16'd0;
            bank111[i] <= 16'd0;
            bank112[i] <= 16'd0;
            bank113[i] <= 16'd0;
            bank114[i] <= 16'd0;
            bank115[i] <= 16'd0;
            bank116[i] <= 16'd0;
            bank117[i] <= 16'd0;
            bank118[i] <= 16'd0;
            bank119[i] <= 16'd0;
            bank120[i] <= 16'd0;
            bank121[i] <= 16'd0;
            bank122[i] <= 16'd0;
            bank123[i] <= 16'd0;
            bank124[i] <= 16'd0;
            bank125[i] <= 16'd0;
            bank126[i] <= 16'd0;
            bank127[i] <= 16'd0;
            bank128[i] <= 16'd0;
            bank129[i] <= 16'd0;
            bank130[i] <= 16'd0;
            bank131[i] <= 16'd0;
            bank132[i] <= 16'd0;
            bank133[i] <= 16'd0;
            bank134[i] <= 16'd0;
            bank135[i] <= 16'd0;
            bank136[i] <= 16'd0;
            bank137[i] <= 16'd0;
            bank138[i] <= 16'd0;
            bank139[i] <= 16'd0;
            bank140[i] <= 16'd0;
            bank141[i] <= 16'd0;
            bank142[i] <= 16'd0;
            bank143[i] <= 16'd0;
            bank144[i] <= 16'd0;
            bank145[i] <= 16'd0;
            bank146[i] <= 16'd0;
            bank147[i] <= 16'd0;
            bank148[i] <= 16'd0;
            bank149[i] <= 16'd0;
            bank150[i] <= 16'd0;
            bank151[i] <= 16'd0;
            bank152[i] <= 16'd0;
            bank153[i] <= 16'd0;
            bank154[i] <= 16'd0;
            bank155[i] <= 16'd0;
            bank156[i] <= 16'd0;
            bank157[i] <= 16'd0;
            bank158[i] <= 16'd0;
            bank159[i] <= 16'd0;
            bank160[i] <= 16'd0;
            bank161[i] <= 16'd0;
            bank162[i] <= 16'd0;
            bank163[i] <= 16'd0;
            bank164[i] <= 16'd0;
            bank165[i] <= 16'd0;
            bank166[i] <= 16'd0;
            bank167[i] <= 16'd0;
            bank168[i] <= 16'd0;
            bank169[i] <= 16'd0;
            bank170[i] <= 16'd0;
            bank171[i] <= 16'd0;
            bank172[i] <= 16'd0;
            bank173[i] <= 16'd0;
            bank174[i] <= 16'd0;
            bank175[i] <= 16'd0;
            bank176[i] <= 16'd0;
            bank177[i] <= 16'd0;
            bank178[i] <= 16'd0;
            bank179[i] <= 16'd0;
            bank180[i] <= 16'd0;
            bank181[i] <= 16'd0;
            bank182[i] <= 16'd0;
            bank183[i] <= 16'd0;
            bank184[i] <= 16'd0;
            bank185[i] <= 16'd0;
            bank186[i] <= 16'd0;
            bank187[i] <= 16'd0;
            bank188[i] <= 16'd0;
            bank189[i] <= 16'd0;
            bank190[i] <= 16'd0;
            bank191[i] <= 16'd0;
            bank192[i] <= 16'd0;
            bank193[i] <= 16'd0;
            bank194[i] <= 16'd0;
            bank195[i] <= 16'd0;
            bank196[i] <= 16'd0;
            bank197[i] <= 16'd0;
            bank198[i] <= 16'd0;
            bank199[i] <= 16'd0;
            bank200[i] <= 16'd0;
            bank201[i] <= 16'd0;
            bank202[i] <= 16'd0;
            bank203[i] <= 16'd0;
            bank204[i] <= 16'd0;
            bank205[i] <= 16'd0;
            bank206[i] <= 16'd0;
            bank207[i] <= 16'd0;
            bank208[i] <= 16'd0;
            bank209[i] <= 16'd0;
            bank210[i] <= 16'd0;
            bank211[i] <= 16'd0;
            bank212[i] <= 16'd0;
            bank213[i] <= 16'd0;
            bank214[i] <= 16'd0;
            bank215[i] <= 16'd0;
            bank216[i] <= 16'd0;
            bank217[i] <= 16'd0;
            bank218[i] <= 16'd0;
            bank219[i] <= 16'd0;
            bank220[i] <= 16'd0;
            bank221[i] <= 16'd0;
            bank222[i] <= 16'd0;
            bank223[i] <= 16'd0;
            bank224[i] <= 16'd0;
            bank225[i] <= 16'd0;
            bank226[i] <= 16'd0;
            bank227[i] <= 16'd0;
            bank228[i] <= 16'd0;
            bank229[i] <= 16'd0;
            bank230[i] <= 16'd0;
            bank231[i] <= 16'd0;
            bank232[i] <= 16'd0;
            bank233[i] <= 16'd0;
            bank234[i] <= 16'd0;
            bank235[i] <= 16'd0;
            bank236[i] <= 16'd0;
            bank237[i] <= 16'd0;
            bank238[i] <= 16'd0;
            bank239[i] <= 16'd0;
            bank240[i] <= 16'd0;
            bank241[i] <= 16'd0;
            bank242[i] <= 16'd0;
            bank243[i] <= 16'd0;
            bank244[i] <= 16'd0;
            bank245[i] <= 16'd0;
            bank246[i] <= 16'd0;
            bank247[i] <= 16'd0;
            bank248[i] <= 16'd0;
            bank249[i] <= 16'd0;
            bank250[i] <= 16'd0;
            bank251[i] <= 16'd0;
            bank252[i] <= 16'd0;
            bank253[i] <= 16'd0;
            bank254[i] <= 16'd0;
            bank255[i] <= 16'd0;
            bank256[i] <= 16'd0;
        end
    else
        if(wren) begin
            bank1[address] <= datainmem[0];
            bank2[address] <= datainmem[1];
            bank3[address] <= datainmem[2];
            bank4[address] <= datainmem[3];
            bank5[address] <= datainmem[4];
            bank6[address] <= datainmem[5];
            bank7[address] <= datainmem[6];
            bank8[address] <= datainmem[7];
            bank9[address] <= datainmem[8];
            bank10[address] <= datainmem[9];
            bank11[address] <= datainmem[10];
            bank12[address] <= datainmem[11];
            bank13[address] <= datainmem[12];
            bank14[address] <= datainmem[13];
            bank15[address] <= datainmem[14];
            bank16[address] <= datainmem[15];
            bank17[address] <= datainmem[16];
            bank18[address] <= datainmem[17];
            bank19[address] <= datainmem[18];
            bank20[address] <= datainmem[19];
            bank21[address] <= datainmem[20];
            bank22[address] <= datainmem[21];
            bank23[address] <= datainmem[22];
            bank24[address] <= datainmem[23];
            bank25[address] <= datainmem[24];
            bank26[address] <= datainmem[25];
            bank27[address] <= datainmem[26];
            bank28[address] <= datainmem[27];
            bank29[address] <= datainmem[28];
            bank30[address] <= datainmem[29];
            bank31[address] <= datainmem[30];
            bank32[address] <= datainmem[31];
            bank33[address] <= datainmem[32];
            bank34[address] <= datainmem[33];
            bank35[address] <= datainmem[34];
            bank36[address] <= datainmem[35];
            bank37[address] <= datainmem[36];
            bank38[address] <= datainmem[37];
            bank39[address] <= datainmem[38];
            bank40[address] <= datainmem[39];
            bank41[address] <= datainmem[40];
            bank42[address] <= datainmem[41];
            bank43[address] <= datainmem[42];
            bank44[address] <= datainmem[43];
            bank45[address] <= datainmem[44];
            bank46[address] <= datainmem[45];
            bank47[address] <= datainmem[46];
            bank48[address] <= datainmem[47];
            bank49[address] <= datainmem[48];
            bank50[address] <= datainmem[49];
            bank51[address] <= datainmem[50];
            bank52[address] <= datainmem[51];
            bank53[address] <= datainmem[52];
            bank54[address] <= datainmem[53];
            bank55[address] <= datainmem[54];
            bank56[address] <= datainmem[55];
            bank57[address] <= datainmem[56];
            bank58[address] <= datainmem[57];
            bank59[address] <= datainmem[58];
            bank60[address] <= datainmem[59];
            bank61[address] <= datainmem[60];
            bank62[address] <= datainmem[61];
            bank63[address] <= datainmem[62];
            bank64[address] <= datainmem[63];
            bank65[address] <= datainmem[64];
            bank66[address] <= datainmem[65];
            bank67[address] <= datainmem[66];
            bank68[address] <= datainmem[67];
            bank69[address] <= datainmem[68];
            bank70[address] <= datainmem[69];
            bank71[address] <= datainmem[70];
            bank72[address] <= datainmem[71];
            bank73[address] <= datainmem[72];
            bank74[address] <= datainmem[73];
            bank75[address] <= datainmem[74];
            bank76[address] <= datainmem[75];
            bank77[address] <= datainmem[76];
            bank78[address] <= datainmem[77];
            bank79[address] <= datainmem[78];
            bank80[address] <= datainmem[79];
            bank81[address] <= datainmem[80];
            bank82[address] <= datainmem[81];
            bank83[address] <= datainmem[82];
            bank84[address] <= datainmem[83];
            bank85[address] <= datainmem[84];
            bank86[address] <= datainmem[85];
            bank87[address] <= datainmem[86];
            bank88[address] <= datainmem[87];
            bank89[address] <= datainmem[88];
            bank90[address] <= datainmem[89];
            bank91[address] <= datainmem[90];
            bank92[address] <= datainmem[91];
            bank93[address] <= datainmem[92];
            bank94[address] <= datainmem[93];
            bank95[address] <= datainmem[94];
            bank96[address] <= datainmem[95];
            bank97[address] <= datainmem[96];
            bank98[address] <= datainmem[97];
            bank99[address] <= datainmem[98];
            bank100[address] <= datainmem[99];
            bank101[address] <= datainmem[100];
            bank102[address] <= datainmem[101];
            bank103[address] <= datainmem[102];
            bank104[address] <= datainmem[103];
            bank105[address] <= datainmem[104];
            bank106[address] <= datainmem[105];
            bank107[address] <= datainmem[106];
            bank108[address] <= datainmem[107];
            bank109[address] <= datainmem[108];
            bank110[address] <= datainmem[109];
            bank111[address] <= datainmem[110];
            bank112[address] <= datainmem[111];
            bank113[address] <= datainmem[112];
            bank114[address] <= datainmem[113];
            bank115[address] <= datainmem[114];
            bank116[address] <= datainmem[115];
            bank117[address] <= datainmem[116];
            bank118[address] <= datainmem[117];
            bank119[address] <= datainmem[118];
            bank120[address] <= datainmem[119];
            bank121[address] <= datainmem[120];
            bank122[address] <= datainmem[121];
            bank123[address] <= datainmem[122];
            bank124[address] <= datainmem[123];
            bank125[address] <= datainmem[124];
            bank126[address] <= datainmem[125];
            bank127[address] <= datainmem[126];
            bank128[address] <= datainmem[127];
            bank129[address] <= datainmem[128];
            bank130[address] <= datainmem[129];
            bank131[address] <= datainmem[130];
            bank132[address] <= datainmem[131];
            bank133[address] <= datainmem[132];
            bank134[address] <= datainmem[133];
            bank135[address] <= datainmem[134];
            bank136[address] <= datainmem[135];
            bank137[address] <= datainmem[136];
            bank138[address] <= datainmem[137];
            bank139[address] <= datainmem[138];
            bank140[address] <= datainmem[139];
            bank141[address] <= datainmem[140];
            bank142[address] <= datainmem[141];
            bank143[address] <= datainmem[142];
            bank144[address] <= datainmem[143];
            bank145[address] <= datainmem[144];
            bank146[address] <= datainmem[145];
            bank147[address] <= datainmem[146];
            bank148[address] <= datainmem[147];
            bank149[address] <= datainmem[148];
            bank150[address] <= datainmem[149];
            bank151[address] <= datainmem[150];
            bank152[address] <= datainmem[151];
            bank153[address] <= datainmem[152];
            bank154[address] <= datainmem[153];
            bank155[address] <= datainmem[154];
            bank156[address] <= datainmem[155];
            bank157[address] <= datainmem[156];
            bank158[address] <= datainmem[157];
            bank159[address] <= datainmem[158];
            bank160[address] <= datainmem[159];
            bank161[address] <= datainmem[160];
            bank162[address] <= datainmem[161];
            bank163[address] <= datainmem[162];
            bank164[address] <= datainmem[163];
            bank165[address] <= datainmem[164];
            bank166[address] <= datainmem[165];
            bank167[address] <= datainmem[166];
            bank168[address] <= datainmem[167];
            bank169[address] <= datainmem[168];
            bank170[address] <= datainmem[169];
            bank171[address] <= datainmem[170];
            bank172[address] <= datainmem[171];
            bank173[address] <= datainmem[172];
            bank174[address] <= datainmem[173];
            bank175[address] <= datainmem[174];
            bank176[address] <= datainmem[175];
            bank177[address] <= datainmem[176];
            bank178[address] <= datainmem[177];
            bank179[address] <= datainmem[178];
            bank180[address] <= datainmem[179];
            bank181[address] <= datainmem[180];
            bank182[address] <= datainmem[181];
            bank183[address] <= datainmem[182];
            bank184[address] <= datainmem[183];
            bank185[address] <= datainmem[184];
            bank186[address] <= datainmem[185];
            bank187[address] <= datainmem[186];
            bank188[address] <= datainmem[187];
            bank189[address] <= datainmem[188];
            bank190[address] <= datainmem[189];
            bank191[address] <= datainmem[190];
            bank192[address] <= datainmem[191];
            bank193[address] <= datainmem[192];
            bank194[address] <= datainmem[193];
            bank195[address] <= datainmem[194];
            bank196[address] <= datainmem[195];
            bank197[address] <= datainmem[196];
            bank198[address] <= datainmem[197];
            bank199[address] <= datainmem[198];
            bank200[address] <= datainmem[199];
            bank201[address] <= datainmem[200];
            bank202[address] <= datainmem[201];
            bank203[address] <= datainmem[202];
            bank204[address] <= datainmem[203];
            bank205[address] <= datainmem[204];
            bank206[address] <= datainmem[205];
            bank207[address] <= datainmem[206];
            bank208[address] <= datainmem[207];
            bank209[address] <= datainmem[208];
            bank210[address] <= datainmem[209];
            bank211[address] <= datainmem[210];
            bank212[address] <= datainmem[211];
            bank213[address] <= datainmem[212];
            bank214[address] <= datainmem[213];
            bank215[address] <= datainmem[214];
            bank216[address] <= datainmem[215];
            bank217[address] <= datainmem[216];
            bank218[address] <= datainmem[217];
            bank219[address] <= datainmem[218];
            bank220[address] <= datainmem[219];
            bank221[address] <= datainmem[220];
            bank222[address] <= datainmem[221];
            bank223[address] <= datainmem[222];
            bank224[address] <= datainmem[223];
            bank225[address] <= datainmem[224];
            bank226[address] <= datainmem[225];
            bank227[address] <= datainmem[226];
            bank228[address] <= datainmem[227];
            bank229[address] <= datainmem[228];
            bank230[address] <= datainmem[229];
            bank231[address] <= datainmem[230];
            bank232[address] <= datainmem[231];
            bank233[address] <= datainmem[232];
            bank234[address] <= datainmem[233];
            bank235[address] <= datainmem[234];
            bank236[address] <= datainmem[235];
            bank237[address] <= datainmem[236];
            bank238[address] <= datainmem[237];
            bank239[address] <= datainmem[238];
            bank240[address] <= datainmem[239];
            bank241[address] <= datainmem[240];
            bank242[address] <= datainmem[241];
            bank243[address] <= datainmem[242];
            bank244[address] <= datainmem[243];
            bank245[address] <= datainmem[244];
            bank246[address] <= datainmem[245];
            bank247[address] <= datainmem[246];
            bank248[address] <= datainmem[247];
            bank249[address] <= datainmem[248];
            bank250[address] <= datainmem[249];
            bank251[address] <= datainmem[250];
            bank252[address] <= datainmem[251];
            bank253[address] <= datainmem[252];
            bank254[address] <= datainmem[253];
            bank255[address] <= datainmem[254];
            bank256[address] <= datainmem[255];
        end
end
always @(*)
begin
    if (rden) begin
    dataoutmem[0] <= bank1[address2];
    dataoutmem[1] <= bank2[address2];
    dataoutmem[2] <= bank3[address2];
    dataoutmem[3] <= bank4[address2];
    dataoutmem[4] <= bank5[address2];
    dataoutmem[5] <= bank6[address2];
    dataoutmem[6] <= bank7[address2];
    dataoutmem[7] <= bank8[address2];
    dataoutmem[8] <= bank9[address2];
    dataoutmem[9] <= bank10[address2];
    dataoutmem[10] <= bank11[address2];
    dataoutmem[11] <= bank12[address2];
    dataoutmem[12] <= bank13[address2];
    dataoutmem[13] <= bank14[address2];
    dataoutmem[14] <= bank15[address2];
    dataoutmem[15] <= bank16[address2];
    dataoutmem[16] <= bank17[address2];
    dataoutmem[17] <= bank18[address2];
    dataoutmem[18] <= bank19[address2];
    dataoutmem[19] <= bank20[address2];
    dataoutmem[20] <= bank21[address2];
    dataoutmem[21] <= bank22[address2];
    dataoutmem[22] <= bank23[address2];
    dataoutmem[23] <= bank24[address2];
    dataoutmem[24] <= bank25[address2];
    dataoutmem[25] <= bank26[address2];
    dataoutmem[26] <= bank27[address2];
    dataoutmem[27] <= bank28[address2];
    dataoutmem[28] <= bank29[address2];
    dataoutmem[29] <= bank30[address2];
    dataoutmem[30] <= bank31[address2];
    dataoutmem[31] <= bank32[address2];
    dataoutmem[32] <= bank33[address2];
    dataoutmem[33] <= bank34[address2];
    dataoutmem[34] <= bank35[address2];
    dataoutmem[35] <= bank36[address2];
    dataoutmem[36] <= bank37[address2];
    dataoutmem[37] <= bank38[address2];
    dataoutmem[38] <= bank39[address2];
    dataoutmem[39] <= bank40[address2];
    dataoutmem[40] <= bank41[address2];
    dataoutmem[41] <= bank42[address2];
    dataoutmem[42] <= bank43[address2];
    dataoutmem[43] <= bank44[address2];
    dataoutmem[44] <= bank45[address2];
    dataoutmem[45] <= bank46[address2];
    dataoutmem[46] <= bank47[address2];
    dataoutmem[47] <= bank48[address2];
    dataoutmem[48] <= bank49[address2];
    dataoutmem[49] <= bank50[address2];
    dataoutmem[50] <= bank51[address2];
    dataoutmem[51] <= bank52[address2];
    dataoutmem[52] <= bank53[address2];
    dataoutmem[53] <= bank54[address2];
    dataoutmem[54] <= bank55[address2];
    dataoutmem[55] <= bank56[address2];
    dataoutmem[56] <= bank57[address2];
    dataoutmem[57] <= bank58[address2];
    dataoutmem[58] <= bank59[address2];
    dataoutmem[59] <= bank60[address2];
    dataoutmem[60] <= bank61[address2];
    dataoutmem[61] <= bank62[address2];
    dataoutmem[62] <= bank63[address2];
    dataoutmem[63] <= bank64[address2];
    dataoutmem[64] <= bank65[address2];
    dataoutmem[65] <= bank66[address2];
    dataoutmem[66] <= bank67[address2];
    dataoutmem[67] <= bank68[address2];
    dataoutmem[68] <= bank69[address2];
    dataoutmem[69] <= bank70[address2];
    dataoutmem[70] <= bank71[address2];
    dataoutmem[71] <= bank72[address2];
    dataoutmem[72] <= bank73[address2];
    dataoutmem[73] <= bank74[address2];
    dataoutmem[74] <= bank75[address2];
    dataoutmem[75] <= bank76[address2];
    dataoutmem[76] <= bank77[address2];
    dataoutmem[77] <= bank78[address2];
    dataoutmem[78] <= bank79[address2];
    dataoutmem[79] <= bank80[address2];
    dataoutmem[80] <= bank81[address2];
    dataoutmem[81] <= bank82[address2];
    dataoutmem[82] <= bank83[address2];
    dataoutmem[83] <= bank84[address2];
    dataoutmem[84] <= bank85[address2];
    dataoutmem[85] <= bank86[address2];
    dataoutmem[86] <= bank87[address2];
    dataoutmem[87] <= bank88[address2];
    dataoutmem[88] <= bank89[address2];
    dataoutmem[89] <= bank90[address2];
    dataoutmem[90] <= bank91[address2];
    dataoutmem[91] <= bank92[address2];
    dataoutmem[92] <= bank93[address2];
    dataoutmem[93] <= bank94[address2];
    dataoutmem[94] <= bank95[address2];
    dataoutmem[95] <= bank96[address2];
    dataoutmem[96] <= bank97[address2];
    dataoutmem[97] <= bank98[address2];
    dataoutmem[98] <= bank99[address2];
    dataoutmem[99] <= bank100[address2];
    dataoutmem[100] <= bank101[address2];
    dataoutmem[101] <= bank102[address2];
    dataoutmem[102] <= bank103[address2];
    dataoutmem[103] <= bank104[address2];
    dataoutmem[104] <= bank105[address2];
    dataoutmem[105] <= bank106[address2];
    dataoutmem[106] <= bank107[address2];
    dataoutmem[107] <= bank108[address2];
    dataoutmem[108] <= bank109[address2];
    dataoutmem[109] <= bank110[address2];
    dataoutmem[110] <= bank111[address2];
    dataoutmem[111] <= bank112[address2];
    dataoutmem[112] <= bank113[address2];
    dataoutmem[113] <= bank114[address2];
    dataoutmem[114] <= bank115[address2];
    dataoutmem[115] <= bank116[address2];
    dataoutmem[116] <= bank117[address2];
    dataoutmem[117] <= bank118[address2];
    dataoutmem[118] <= bank119[address2];
    dataoutmem[119] <= bank120[address2];
    dataoutmem[120] <= bank121[address2];
    dataoutmem[121] <= bank122[address2];
    dataoutmem[122] <= bank123[address2];
    dataoutmem[123] <= bank124[address2];
    dataoutmem[124] <= bank125[address2];
    dataoutmem[125] <= bank126[address2];
    dataoutmem[126] <= bank127[address2];
    dataoutmem[127] <= bank128[address2];
    dataoutmem[128] <= bank129[address2];
    dataoutmem[129] <= bank130[address2];
    dataoutmem[130] <= bank131[address2];
    dataoutmem[131] <= bank132[address2];
    dataoutmem[132] <= bank133[address2];
    dataoutmem[133] <= bank134[address2];
    dataoutmem[134] <= bank135[address2];
    dataoutmem[135] <= bank136[address2];
    dataoutmem[136] <= bank137[address2];
    dataoutmem[137] <= bank138[address2];
    dataoutmem[138] <= bank139[address2];
    dataoutmem[139] <= bank140[address2];
    dataoutmem[140] <= bank141[address2];
    dataoutmem[141] <= bank142[address2];
    dataoutmem[142] <= bank143[address2];
    dataoutmem[143] <= bank144[address2];
    dataoutmem[144] <= bank145[address2];
    dataoutmem[145] <= bank146[address2];
    dataoutmem[146] <= bank147[address2];
    dataoutmem[147] <= bank148[address2];
    dataoutmem[148] <= bank149[address2];
    dataoutmem[149] <= bank150[address2];
    dataoutmem[150] <= bank151[address2];
    dataoutmem[151] <= bank152[address2];
    dataoutmem[152] <= bank153[address2];
    dataoutmem[153] <= bank154[address2];
    dataoutmem[154] <= bank155[address2];
    dataoutmem[155] <= bank156[address2];
    dataoutmem[156] <= bank157[address2];
    dataoutmem[157] <= bank158[address2];
    dataoutmem[158] <= bank159[address2];
    dataoutmem[159] <= bank160[address2];
    dataoutmem[160] <= bank161[address2];
    dataoutmem[161] <= bank162[address2];
    dataoutmem[162] <= bank163[address2];
    dataoutmem[163] <= bank164[address2];
    dataoutmem[164] <= bank165[address2];
    dataoutmem[165] <= bank166[address2];
    dataoutmem[166] <= bank167[address2];
    dataoutmem[167] <= bank168[address2];
    dataoutmem[168] <= bank169[address2];
    dataoutmem[169] <= bank170[address2];
    dataoutmem[170] <= bank171[address2];
    dataoutmem[171] <= bank172[address2];
    dataoutmem[172] <= bank173[address2];
    dataoutmem[173] <= bank174[address2];
    dataoutmem[174] <= bank175[address2];
    dataoutmem[175] <= bank176[address2];
    dataoutmem[176] <= bank177[address2];
    dataoutmem[177] <= bank178[address2];
    dataoutmem[178] <= bank179[address2];
    dataoutmem[179] <= bank180[address2];
    dataoutmem[180] <= bank181[address2];
    dataoutmem[181] <= bank182[address2];
    dataoutmem[182] <= bank183[address2];
    dataoutmem[183] <= bank184[address2];
    dataoutmem[184] <= bank185[address2];
    dataoutmem[185] <= bank186[address2];
    dataoutmem[186] <= bank187[address2];
    dataoutmem[187] <= bank188[address2];
    dataoutmem[188] <= bank189[address2];
    dataoutmem[189] <= bank190[address2];
    dataoutmem[190] <= bank191[address2];
    dataoutmem[191] <= bank192[address2];
    dataoutmem[192] <= bank193[address2];
    dataoutmem[193] <= bank194[address2];
    dataoutmem[194] <= bank195[address2];
    dataoutmem[195] <= bank196[address2];
    dataoutmem[196] <= bank197[address2];
    dataoutmem[197] <= bank198[address2];
    dataoutmem[198] <= bank199[address2];
    dataoutmem[199] <= bank200[address2];
    dataoutmem[200] <= bank201[address2];
    dataoutmem[201] <= bank202[address2];
    dataoutmem[202] <= bank203[address2];
    dataoutmem[203] <= bank204[address2];
    dataoutmem[204] <= bank205[address2];
    dataoutmem[205] <= bank206[address2];
    dataoutmem[206] <= bank207[address2];
    dataoutmem[207] <= bank208[address2];
    dataoutmem[208] <= bank209[address2];
    dataoutmem[209] <= bank210[address2];
    dataoutmem[210] <= bank211[address2];
    dataoutmem[211] <= bank212[address2];
    dataoutmem[212] <= bank213[address2];
    dataoutmem[213] <= bank214[address2];
    dataoutmem[214] <= bank215[address2];
    dataoutmem[215] <= bank216[address2];
    dataoutmem[216] <= bank217[address2];
    dataoutmem[217] <= bank218[address2];
    dataoutmem[218] <= bank219[address2];
    dataoutmem[219] <= bank220[address2];
    dataoutmem[220] <= bank221[address2];
    dataoutmem[221] <= bank222[address2];
    dataoutmem[222] <= bank223[address2];
    dataoutmem[223] <= bank224[address2];
    dataoutmem[224] <= bank225[address2];
    dataoutmem[225] <= bank226[address2];
    dataoutmem[226] <= bank227[address2];
    dataoutmem[227] <= bank228[address2];
    dataoutmem[228] <= bank229[address2];
    dataoutmem[229] <= bank230[address2];
    dataoutmem[230] <= bank231[address2];
    dataoutmem[231] <= bank232[address2];
    dataoutmem[232] <= bank233[address2];
    dataoutmem[233] <= bank234[address2];
    dataoutmem[234] <= bank235[address2];
    dataoutmem[235] <= bank236[address2];
    dataoutmem[236] <= bank237[address2];
    dataoutmem[237] <= bank238[address2];
    dataoutmem[238] <= bank239[address2];
    dataoutmem[239] <= bank240[address2];
    dataoutmem[240] <= bank241[address2];
    dataoutmem[241] <= bank242[address2];
    dataoutmem[242] <= bank243[address2];
    dataoutmem[243] <= bank244[address2];
    dataoutmem[244] <= bank245[address2];
    dataoutmem[245] <= bank246[address2];
    dataoutmem[246] <= bank247[address2];
    dataoutmem[247] <= bank248[address2];
    dataoutmem[248] <= bank249[address2];
    dataoutmem[249] <= bank250[address2];
    dataoutmem[250] <= bank251[address2];
    dataoutmem[251] <= bank252[address2];
    dataoutmem[252] <= bank253[address2];
    dataoutmem[253] <= bank254[address2];
    dataoutmem[254] <= bank255[address2];
    dataoutmem[255] <= bank256[address2];
    end
end
always @(*)
begin
for (i=0; i<256; i=i+1)
    dataout[i*16+:16]<=dataoutmem[i];
end
endmodule