module conv1banks(clk,rst, wren, rden, address, address2, datain, dataout);
input clk, rst;
reg [15:0] bank1 [0:111*111-1];
reg [15:0] bank2 [0:111*111-1];
reg [15:0] bank3 [0:111*111-1];
reg [15:0] bank4 [0:111*111-1];
reg [15:0] bank5 [0:111*111-1];
reg [15:0] bank6 [0:111*111-1];
reg [15:0] bank7 [0:111*111-1];
reg [15:0] bank8 [0:111*111-1];
reg [15:0] bank9 [0:111*111-1];
reg [15:0] bank10 [0:111*111-1];
reg [15:0] bank11 [0:111*111-1];
reg [15:0] bank12 [0:111*111-1];
reg [15:0] bank13 [0:111*111-1];
reg [15:0] bank14 [0:111*111-1];
reg [15:0] bank15 [0:111*111-1];
reg [15:0] bank16 [0:111*111-1];
reg [15:0] bank17 [0:111*111-1];
reg [15:0] bank18 [0:111*111-1];
reg [15:0] bank19 [0:111*111-1];
reg [15:0] bank20 [0:111*111-1];
reg [15:0] bank21 [0:111*111-1];
reg [15:0] bank22 [0:111*111-1];
reg [15:0] bank23 [0:111*111-1];
reg [15:0] bank24 [0:111*111-1];
reg [15:0] bank25 [0:111*111-1];
reg [15:0] bank26 [0:111*111-1];
reg [15:0] bank27 [0:111*111-1];
reg [15:0] bank28 [0:111*111-1];
reg [15:0] bank29 [0:111*111-1];
reg [15:0] bank30 [0:111*111-1];
reg [15:0] bank31 [0:111*111-1];
reg [15:0] bank32 [0:111*111-1];
reg [15:0] bank33 [0:111*111-1];
reg [15:0] bank34 [0:111*111-1];
reg [15:0] bank35 [0:111*111-1];
reg [15:0] bank36 [0:111*111-1];
reg [15:0] bank37 [0:111*111-1];
reg [15:0] bank38 [0:111*111-1];
reg [15:0] bank39 [0:111*111-1];
reg [15:0] bank40 [0:111*111-1];
reg [15:0] bank41 [0:111*111-1];
reg [15:0] bank42 [0:111*111-1];
reg [15:0] bank43 [0:111*111-1];
reg [15:0] bank44 [0:111*111-1];
reg [15:0] bank45 [0:111*111-1];
reg [15:0] bank46 [0:111*111-1];
reg [15:0] bank47 [0:111*111-1];
reg [15:0] bank48 [0:111*111-1];
reg [15:0] bank49 [0:111*111-1];
reg [15:0] bank50 [0:111*111-1];
reg [15:0] bank51 [0:111*111-1];
reg [15:0] bank52 [0:111*111-1];
reg [15:0] bank53 [0:111*111-1];
reg [15:0] bank54 [0:111*111-1];
reg [15:0] bank55 [0:111*111-1];
reg [15:0] bank56 [0:111*111-1];
reg [15:0] bank57 [0:111*111-1];
reg [15:0] bank58 [0:111*111-1];
reg [15:0] bank59 [0:111*111-1];
reg [15:0] bank60 [0:111*111-1];
reg [15:0] bank61 [0:111*111-1];
reg [15:0] bank62 [0:111*111-1];
reg [15:0] bank63 [0:111*111-1];
reg [15:0] bank64 [0:111*111-1];


input rden;
input wren;
input [32-1:0] address;
input [32-1:0] address2;
input [16*64-1:0] datain;
reg [15:0] datainmem[0:63];
output reg [16*64-1:0] dataout;
reg [15:0] dataoutmem[0:63];
integer i;
always @(*)
begin
for (i=0; i<64; i=i+1)
    datainmem[i]<=datain[i*16+:16];
end
always @(posedge clk)
begin
    if(rst)
        for (i=0; i<111*111;i=i+1) begin
            bank1[i] <= 16'd0;
            bank2[i] <= 16'd0;
            bank3[i] <= 16'd0;
            bank4[i] <= 16'd0;
            bank5[i] <= 16'd0;
            bank6[i] <= 16'd0;
            bank7[i] <= 16'd0;
            bank8[i] <= 16'd0;
            bank9[i] <= 16'd0;
            bank10[i] <= 16'd0;
            bank11[i] <= 16'd0;
            bank12[i] <= 16'd0;
            bank13[i] <= 16'd0;
            bank14[i] <= 16'd0;
            bank15[i] <= 16'd0;
            bank16[i] <= 16'd0;
            bank17[i] <= 16'd0;
            bank18[i] <= 16'd0;
            bank19[i] <= 16'd0;
            bank20[i] <= 16'd0;
            bank21[i] <= 16'd0;
            bank22[i] <= 16'd0;
            bank23[i] <= 16'd0;
            bank24[i] <= 16'd0;
            bank25[i] <= 16'd0;
            bank26[i] <= 16'd0;
            bank27[i] <= 16'd0;
            bank28[i] <= 16'd0;
            bank29[i] <= 16'd0;
            bank30[i] <= 16'd0;
            bank31[i] <= 16'd0;
            bank32[i] <= 16'd0;
            bank33[i] <= 16'd0;
            bank34[i] <= 16'd0;
            bank35[i] <= 16'd0;
            bank36[i] <= 16'd0;
            bank37[i] <= 16'd0;
            bank38[i] <= 16'd0;
            bank39[i] <= 16'd0;
            bank40[i] <= 16'd0;
            bank41[i] <= 16'd0;
            bank42[i] <= 16'd0;
            bank43[i] <= 16'd0;
            bank44[i] <= 16'd0;
            bank45[i] <= 16'd0;
            bank46[i] <= 16'd0;
            bank47[i] <= 16'd0;
            bank48[i] <= 16'd0;
            bank49[i] <= 16'd0;
            bank50[i] <= 16'd0;
            bank51[i] <= 16'd0;
            bank52[i] <= 16'd0;
            bank53[i] <= 16'd0;
            bank54[i] <= 16'd0;
            bank55[i] <= 16'd0;
            bank56[i] <= 16'd0;
            bank57[i] <= 16'd0;
            bank58[i] <= 16'd0;
            bank59[i] <= 16'd0;
            bank60[i] <= 16'd0;
            bank61[i] <= 16'd0;
            bank62[i] <= 16'd0;
            bank63[i] <= 16'd0;
            bank64[i] <= 16'd0;
        end
    else
        if(wren) begin
            bank1[address] <= datainmem[0];
            bank2[address] <= datainmem[1];
            bank3[address] <= datainmem[2];
            bank4[address] <= datainmem[3];
            bank5[address] <= datainmem[4];
            bank6[address] <= datainmem[5];
            bank7[address] <= datainmem[6];
            bank8[address] <= datainmem[7];
            bank9[address] <= datainmem[8];
            bank10[address] <= datainmem[9];
            bank11[address] <= datainmem[10];
            bank12[address] <= datainmem[11];
            bank13[address] <= datainmem[12];
            bank14[address] <= datainmem[13];
            bank15[address] <= datainmem[14];
            bank16[address] <= datainmem[15];
            bank17[address] <= datainmem[16];
            bank18[address] <= datainmem[17];
            bank19[address] <= datainmem[18];
            bank20[address] <= datainmem[19];
            bank21[address] <= datainmem[20];
            bank22[address] <= datainmem[21];
            bank23[address] <= datainmem[22];
            bank24[address] <= datainmem[23];
            bank25[address] <= datainmem[24];
            bank26[address] <= datainmem[25];
            bank27[address] <= datainmem[26];
            bank28[address] <= datainmem[27];
            bank29[address] <= datainmem[28];
            bank30[address] <= datainmem[29];
            bank31[address] <= datainmem[30];
            bank32[address] <= datainmem[31];
            bank33[address] <= datainmem[32];
            bank34[address] <= datainmem[33];
            bank35[address] <= datainmem[34];
            bank36[address] <= datainmem[35];
            bank37[address] <= datainmem[36];
            bank38[address] <= datainmem[37];
            bank39[address] <= datainmem[38];
            bank40[address] <= datainmem[39];
            bank41[address] <= datainmem[40];
            bank42[address] <= datainmem[41];
            bank43[address] <= datainmem[42];
            bank44[address] <= datainmem[43];
            bank45[address] <= datainmem[44];
            bank46[address] <= datainmem[45];
            bank47[address] <= datainmem[46];
            bank48[address] <= datainmem[47];
            bank49[address] <= datainmem[48];
            bank50[address] <= datainmem[49];
            bank51[address] <= datainmem[50];
            bank52[address] <= datainmem[51];
            bank53[address] <= datainmem[52];
            bank54[address] <= datainmem[53];
            bank55[address] <= datainmem[54];
            bank56[address] <= datainmem[55];
            bank57[address] <= datainmem[56];
            bank58[address] <= datainmem[57];
            bank59[address] <= datainmem[58];
            bank60[address] <= datainmem[59];
            bank61[address] <= datainmem[60];
            bank62[address] <= datainmem[61];
            bank63[address] <= datainmem[62];
            bank64[address] <= datainmem[63];
        end
end
always @(*)
begin
if (rden) begin
    dataoutmem[0] <= bank1[address2];
    dataoutmem[1] <= bank2[address2];
    dataoutmem[2] <= bank3[address2];
    dataoutmem[3] <= bank4[address2];
    dataoutmem[4] <= bank5[address2];
    dataoutmem[5] <= bank6[address2];
    dataoutmem[6] <= bank7[address2];
    dataoutmem[7] <= bank8[address2];
    dataoutmem[8] <= bank9[address2];
    dataoutmem[9] <= bank10[address2];
    dataoutmem[10] <= bank11[address2];
    dataoutmem[11] <= bank12[address2];
    dataoutmem[12] <= bank13[address2];
    dataoutmem[13] <= bank14[address2];
    dataoutmem[14] <= bank15[address2];
    dataoutmem[15] <= bank16[address2];
    dataoutmem[16] <= bank17[address2];
    dataoutmem[17] <= bank18[address2];
    dataoutmem[18] <= bank19[address2];
    dataoutmem[19] <= bank20[address2];
    dataoutmem[20] <= bank21[address2];
    dataoutmem[21] <= bank22[address2];
    dataoutmem[22] <= bank23[address2];
    dataoutmem[23] <= bank24[address2];
    dataoutmem[24] <= bank25[address2];
    dataoutmem[25] <= bank26[address2];
    dataoutmem[26] <= bank27[address2];
    dataoutmem[27] <= bank28[address2];
    dataoutmem[28] <= bank29[address2];
    dataoutmem[29] <= bank30[address2];
    dataoutmem[30] <= bank31[address2];
    dataoutmem[31] <= bank32[address2];
    dataoutmem[32] <= bank33[address2];
    dataoutmem[33] <= bank34[address2];
    dataoutmem[34] <= bank35[address2];
    dataoutmem[35] <= bank36[address2];
    dataoutmem[36] <= bank37[address2];
    dataoutmem[37] <= bank38[address2];
    dataoutmem[38] <= bank39[address2];
    dataoutmem[39] <= bank40[address2];
    dataoutmem[40] <= bank41[address2];
    dataoutmem[41] <= bank42[address2];
    dataoutmem[42] <= bank43[address2];
    dataoutmem[43] <= bank44[address2];
    dataoutmem[44] <= bank45[address2];
    dataoutmem[45] <= bank46[address2];
    dataoutmem[46] <= bank47[address2];
    dataoutmem[47] <= bank48[address2];
    dataoutmem[48] <= bank49[address2];
    dataoutmem[49] <= bank50[address2];
    dataoutmem[50] <= bank51[address2];
    dataoutmem[51] <= bank52[address2];
    dataoutmem[52] <= bank53[address2];
    dataoutmem[53] <= bank54[address2];
    dataoutmem[54] <= bank55[address2];
    dataoutmem[55] <= bank56[address2];
    dataoutmem[56] <= bank57[address2];
    dataoutmem[57] <= bank58[address2];
    dataoutmem[58] <= bank59[address2];
    dataoutmem[59] <= bank60[address2];
    dataoutmem[60] <= bank61[address2];
    dataoutmem[61] <= bank62[address2];
    dataoutmem[62] <= bank63[address2];
    dataoutmem[63] <= bank64[address2];
end
end
always @(*)
begin
for (i=0; i<64; i=i+1)
    dataout[i*16+:16]<=dataoutmem[i];
end
endmodule