module maxpool2d(clk, rst, i_data_valid, pooladdr, inp,maxpoolout,maxpoolvalid);
input [64*16-1:0] inp;
reg [15:0] inpmem [0:64-1];
output reg [64*16-1:0] maxpoolout;
wire [15:0] maxpooloutmem [0:64-1];
output maxpoolvalid;
wire [63:0] maxpooloutvalid;
output [31:0] pooladdr;
input clk, rst, i_data_valid;
integer i;
always @(*)
begin
for (i=0; i<64; i=i+1)
    inpmem[i]<=inp[i*16+:16];
end
maxpool2d3x3 maxpool (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[0]),.address(pooladdr),.output_im(maxpooloutmem[0]),.o_max_data_valid(maxpooloutvalid[0]));
maxpool2d3x3 maxpool1 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[1]),.address(pooladdr),.output_im(maxpooloutmem[1]),.o_max_data_valid(maxpooloutvalid[1]));
maxpool2d3x3 maxpool2 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[2]),.address(pooladdr),.output_im(maxpooloutmem[2]),.o_max_data_valid(maxpooloutvalid[2]));
maxpool2d3x3 maxpool3 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[3]),.address(pooladdr),.output_im(maxpooloutmem[3]),.o_max_data_valid(maxpooloutvalid[3]));
maxpool2d3x3 maxpool4 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[4]),.address(pooladdr),.output_im(maxpooloutmem[4]),.o_max_data_valid(maxpooloutvalid[4]));
maxpool2d3x3 maxpool5 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[5]),.address(pooladdr),.output_im(maxpooloutmem[5]),.o_max_data_valid(maxpooloutvalid[5]));
maxpool2d3x3 maxpool6 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[6]),.address(pooladdr),.output_im(maxpooloutmem[6]),.o_max_data_valid(maxpooloutvalid[6]));
maxpool2d3x3 maxpool7 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[7]),.address(pooladdr),.output_im(maxpooloutmem[7]),.o_max_data_valid(maxpooloutvalid[7]));
maxpool2d3x3 maxpool8 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[8]),.address(pooladdr),.output_im(maxpooloutmem[8]),.o_max_data_valid(maxpooloutvalid[8]));
maxpool2d3x3 maxpool9 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[9]),.address(pooladdr),.output_im(maxpooloutmem[9]),.o_max_data_valid(maxpooloutvalid[9]));
maxpool2d3x3 maxpool10 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[10]),.address(pooladdr),.output_im(maxpooloutmem[10]),.o_max_data_valid(maxpooloutvalid[10]));
maxpool2d3x3 maxpool11 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[11]),.address(pooladdr),.output_im(maxpooloutmem[11]),.o_max_data_valid(maxpooloutvalid[11]));
maxpool2d3x3 maxpool12 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[12]),.address(pooladdr),.output_im(maxpooloutmem[12]),.o_max_data_valid(maxpooloutvalid[12]));
maxpool2d3x3 maxpool13 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[13]),.address(pooladdr),.output_im(maxpooloutmem[13]),.o_max_data_valid(maxpooloutvalid[13]));
maxpool2d3x3 maxpool14 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[14]),.address(pooladdr),.output_im(maxpooloutmem[14]),.o_max_data_valid(maxpooloutvalid[14]));
maxpool2d3x3 maxpool15 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[15]),.address(pooladdr),.output_im(maxpooloutmem[15]),.o_max_data_valid(maxpooloutvalid[15]));
maxpool2d3x3 maxpool16 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[16]),.address(pooladdr),.output_im(maxpooloutmem[16]),.o_max_data_valid(maxpooloutvalid[16]));
maxpool2d3x3 maxpool17 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[17]),.address(pooladdr),.output_im(maxpooloutmem[17]),.o_max_data_valid(maxpooloutvalid[17]));
maxpool2d3x3 maxpool18 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[18]),.address(pooladdr),.output_im(maxpooloutmem[18]),.o_max_data_valid(maxpooloutvalid[18]));
maxpool2d3x3 maxpool19 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[19]),.address(pooladdr),.output_im(maxpooloutmem[19]),.o_max_data_valid(maxpooloutvalid[19]));
maxpool2d3x3 maxpool20 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[20]),.address(pooladdr),.output_im(maxpooloutmem[20]),.o_max_data_valid(maxpooloutvalid[20]));
maxpool2d3x3 maxpool21 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[21]),.address(pooladdr),.output_im(maxpooloutmem[21]),.o_max_data_valid(maxpooloutvalid[21]));
maxpool2d3x3 maxpool22 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[22]),.address(pooladdr),.output_im(maxpooloutmem[22]),.o_max_data_valid(maxpooloutvalid[22]));
maxpool2d3x3 maxpool23 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[23]),.address(pooladdr),.output_im(maxpooloutmem[23]),.o_max_data_valid(maxpooloutvalid[23]));
maxpool2d3x3 maxpool24 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[24]),.address(pooladdr),.output_im(maxpooloutmem[24]),.o_max_data_valid(maxpooloutvalid[24]));
maxpool2d3x3 maxpool25 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[25]),.address(pooladdr),.output_im(maxpooloutmem[25]),.o_max_data_valid(maxpooloutvalid[25]));
maxpool2d3x3 maxpool26 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[26]),.address(pooladdr),.output_im(maxpooloutmem[26]),.o_max_data_valid(maxpooloutvalid[26]));
maxpool2d3x3 maxpool27 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[27]),.address(pooladdr),.output_im(maxpooloutmem[27]),.o_max_data_valid(maxpooloutvalid[27]));
maxpool2d3x3 maxpool28 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[28]),.address(pooladdr),.output_im(maxpooloutmem[28]),.o_max_data_valid(maxpooloutvalid[28]));
maxpool2d3x3 maxpool29 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[29]),.address(pooladdr),.output_im(maxpooloutmem[29]),.o_max_data_valid(maxpooloutvalid[29]));
maxpool2d3x3 maxpool30 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[30]),.address(pooladdr),.output_im(maxpooloutmem[30]),.o_max_data_valid(maxpooloutvalid[30]));
maxpool2d3x3 maxpool31 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[31]),.address(pooladdr),.output_im(maxpooloutmem[31]),.o_max_data_valid(maxpooloutvalid[31]));
maxpool2d3x3 maxpool32 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[32]),.address(pooladdr),.output_im(maxpooloutmem[32]),.o_max_data_valid(maxpooloutvalid[32]));
maxpool2d3x3 maxpool33 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[33]),.address(pooladdr),.output_im(maxpooloutmem[33]),.o_max_data_valid(maxpooloutvalid[33]));
maxpool2d3x3 maxpool34 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[34]),.address(pooladdr),.output_im(maxpooloutmem[34]),.o_max_data_valid(maxpooloutvalid[34]));
maxpool2d3x3 maxpool35 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[35]),.address(pooladdr),.output_im(maxpooloutmem[35]),.o_max_data_valid(maxpooloutvalid[35]));
maxpool2d3x3 maxpool36 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[36]),.address(pooladdr),.output_im(maxpooloutmem[36]),.o_max_data_valid(maxpooloutvalid[36]));
maxpool2d3x3 maxpool37 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[37]),.address(pooladdr),.output_im(maxpooloutmem[37]),.o_max_data_valid(maxpooloutvalid[37]));
maxpool2d3x3 maxpool38 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[38]),.address(pooladdr),.output_im(maxpooloutmem[38]),.o_max_data_valid(maxpooloutvalid[38]));
maxpool2d3x3 maxpool39 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[39]),.address(pooladdr),.output_im(maxpooloutmem[39]),.o_max_data_valid(maxpooloutvalid[39]));
maxpool2d3x3 maxpool40 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[40]),.address(pooladdr),.output_im(maxpooloutmem[40]),.o_max_data_valid(maxpooloutvalid[40]));
maxpool2d3x3 maxpool41 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[41]),.address(pooladdr),.output_im(maxpooloutmem[41]),.o_max_data_valid(maxpooloutvalid[41]));
maxpool2d3x3 maxpool42 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[42]),.address(pooladdr),.output_im(maxpooloutmem[42]),.o_max_data_valid(maxpooloutvalid[42]));
maxpool2d3x3 maxpool43 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[43]),.address(pooladdr),.output_im(maxpooloutmem[43]),.o_max_data_valid(maxpooloutvalid[43]));
maxpool2d3x3 maxpool44 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[44]),.address(pooladdr),.output_im(maxpooloutmem[44]),.o_max_data_valid(maxpooloutvalid[44]));
maxpool2d3x3 maxpool45 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[45]),.address(pooladdr),.output_im(maxpooloutmem[45]),.o_max_data_valid(maxpooloutvalid[45]));
maxpool2d3x3 maxpool46 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[46]),.address(pooladdr),.output_im(maxpooloutmem[46]),.o_max_data_valid(maxpooloutvalid[46]));
maxpool2d3x3 maxpool47 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[47]),.address(pooladdr),.output_im(maxpooloutmem[47]),.o_max_data_valid(maxpooloutvalid[47]));
maxpool2d3x3 maxpool48 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[48]),.address(pooladdr),.output_im(maxpooloutmem[48]),.o_max_data_valid(maxpooloutvalid[48]));
maxpool2d3x3 maxpool49 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[49]),.address(pooladdr),.output_im(maxpooloutmem[49]),.o_max_data_valid(maxpooloutvalid[49]));
maxpool2d3x3 maxpool50 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[50]),.address(pooladdr),.output_im(maxpooloutmem[50]),.o_max_data_valid(maxpooloutvalid[50]));
maxpool2d3x3 maxpool51 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[51]),.address(pooladdr),.output_im(maxpooloutmem[51]),.o_max_data_valid(maxpooloutvalid[51]));
maxpool2d3x3 maxpool52 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[52]),.address(pooladdr),.output_im(maxpooloutmem[52]),.o_max_data_valid(maxpooloutvalid[52]));
maxpool2d3x3 maxpool53 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[53]),.address(pooladdr),.output_im(maxpooloutmem[53]),.o_max_data_valid(maxpooloutvalid[53]));
maxpool2d3x3 maxpool54 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[54]),.address(pooladdr),.output_im(maxpooloutmem[54]),.o_max_data_valid(maxpooloutvalid[54]));
maxpool2d3x3 maxpool55 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[55]),.address(pooladdr),.output_im(maxpooloutmem[55]),.o_max_data_valid(maxpooloutvalid[55]));
maxpool2d3x3 maxpool56 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[56]),.address(pooladdr),.output_im(maxpooloutmem[56]),.o_max_data_valid(maxpooloutvalid[56]));
maxpool2d3x3 maxpool57 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[57]),.address(pooladdr),.output_im(maxpooloutmem[57]),.o_max_data_valid(maxpooloutvalid[57]));
maxpool2d3x3 maxpool58 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[58]),.address(pooladdr),.output_im(maxpooloutmem[58]),.o_max_data_valid(maxpooloutvalid[58]));
maxpool2d3x3 maxpool59 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[59]),.address(pooladdr),.output_im(maxpooloutmem[59]),.o_max_data_valid(maxpooloutvalid[59]));
maxpool2d3x3 maxpool60 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[60]),.address(pooladdr),.output_im(maxpooloutmem[60]),.o_max_data_valid(maxpooloutvalid[60]));
maxpool2d3x3 maxpool61 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[61]),.address(pooladdr),.output_im(maxpooloutmem[61]),.o_max_data_valid(maxpooloutvalid[61]));
maxpool2d3x3 maxpool62 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[62]),.address(pooladdr),.output_im(maxpooloutmem[62]),.o_max_data_valid(maxpooloutvalid[62]));
maxpool2d3x3 maxpool63 (.clk(clk),.rst(rst),.i_data_valid(i_data_valid),.datain(inpmem[63]),.address(pooladdr),.output_im(maxpooloutmem[63]),.o_max_data_valid(maxpooloutvalid[63]));

assign maxpoolvalid=|maxpooloutvalid;
always @(*)
begin
for (i=0; i<64; i=i+1)
    maxpoolout[i*16+:16]<=maxpooloutmem[i];
end
endmodule